	module clk_div (WIDTH, N, clk,reset, slow_clk);
  
	input WIDTH = 3, // Width of the register required
	input N = 6// We will divide by 12 for example in this case
	input clk;
	input reset;
	output slow_clk;
	 
	reg [WIDTH-1:0] r_reg;
	wire [WIDTH-1:0] r_nxt;
	reg clk_track;
	 
	always @(posedge clk or posedge reset)
	 
	begin
	  if (reset)
	     begin
	        r_reg <= 0;
	      clk_track <= 1'b0;
	     end
	 
	  else if (r_nxt == N)
	        begin
	           r_reg <= 0;
	           clk_track <= ~clk_track;
	         end
	 
	  else 
	      r_reg <= r_nxt;
	end
	 
	assign r_nxt = r_reg+1;            
	assign slow_clk = clk_track;
endmodule
