module main();
	input KEY0, KEY1, KEY2, KEY3;
	output [0:9] LEDR;
	seg_disp display();
endmodule
