module seg_disp
(
  input [9:0] SW,
  output [0:6] HEX0, HEX1, HEX2, HEX3,
  output [0:9] LEDR
);
 
endmodule
