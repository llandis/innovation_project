module sequencer(
input pb_seq_up;
input pb_seq_dn;
input slow_clk;
input clk_50;
input reset;

output ROM_addr;
output seq_num;
output LEDS;
);



end
