module sequencer(
input CLK_50,
input reset,
input pb_freq_up,
input pb_freq_dn,

output slow_clk,
output freq_num,
);

endmodule
