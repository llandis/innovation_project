// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 16.0.0 Build 211 04/27/2016 SJ Standard Edition
// Created on Wed Nov  2 11:10:02 2016

// synthesis message_off 10175

`timescale 1ns/1ns

module ROM_state (
    reset_n,clock_n,length[5:0],start[9:0],end_seq[9:0],at_end,first_ram,last_ram,pb_seq_up,pb_seq_dn,reset,
    load,addr[9:0],ram_counter[5:0],at_end_rst,addr_inc,ram_counter_inc,ram_counter_dec);

    input reset_n;
    input clock_n;
    input [5:0] length;
    input [9:0] start;
	input [9:0] end_seq;
	 input at_end;
	 input first_ram;
	 input last_ram;
	 input pb_seq_up;
	 input pb_seq_dn;
	 input reset;
    tri0 reset_n;
    tri0 [5:0] length;
    tri0 [9:0] start;
	tri0 [9:0] end_seq;
	 tri0 at_end;
	 tri0 first_ram;
	 tri0 last_ram;
	 tri0 pb_seq_up;
	 tri0 pb_seq_dn;
	 tri0 reset;
    output load;
    output [9:0] addr;
    output [5:0] ram_counter;
    output at_end_rst;
    output addr_inc;
    output ram_counter_inc;
    output ram_counter_dec;
    reg load;
    reg [9:0] addr;
    reg [5:0] ram_counter;
    reg at_end_rst;
    reg addr_inc;
    reg ram_counter_inc;
    reg ram_counter_dec;
    reg [5:0] fstate;
    reg [5:0] reg_fstate;
    parameter INIT=0,IN_SEQ=1,BOT_SEQ=2,NEXT_SEQ=3,PREV_SEQ=4,LAST_SEQ=5;

    always @(posedge clock_n)
    begin
        if (clock_n) begin
            fstate <= reg_fstate;
        end
    end
	
	always @(posedge clock_n)
	begin
		if(load == 1'b1) begin
			//write logic to reference the correct start number
			//put the start number inside addr
		end
		
		at_end = and(~at_end_rst, end_seq, addr)

    always @(fstate or reset_n or length or start or end_seq or at_end or first_ram or last_ram or pb_seq_up or pb_seq_dn or reset)
    begin
        if (reset) begin
            reg_fstate <= INIT;
            load <= 1'b0;
            addr <= 10'b0000000000;
            ram_counter <= 6'b000000;
            at_end_rst <= 1'b0;
            addr_inc <= 1'b0;
            ram_counter_inc <= 1'b0;
            ram_counter_dec <= 1'b0;
        end
        else begin
            load <= 1'b0;
            addr <= 10'b0000000000;
            ram_counter <= 6'b000000;
            at_end_rst <= 1'b0;
            addr_inc <= 1'b0;
            ram_counter_inc <= 1'b0;
            ram_counter_dec <= 1'b0;
            case (fstate)
                INIT: begin
                    if ((reset == 1'b0))
                        reg_fstate <= IN_SEQ;
                    else if ((reset == 1'b1))
                        reg_fstate <= INIT;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= INIT;

                    at_end_rst <= 1'b0;
                    ram_counter <= 6'b000000;

                    //addr <= start[9:0];

                    load <= 1'b0;
                end
                IN_SEQ: begin
                    if ((pb_seq_dn == 1'b1 && pb_seq_up == 1'b0))
                        reg_fstate <= PREV_SEQ;
                    else if ((pb_seq_up == 1'b1 && pb_seq_dn == 1'b0))
                        reg_fstate <= NEXT_SEQ;
                    else if ((pb_seq_dn == 1'b1 && addr == 10'b00_0000_0000))
                        reg_fstate <= LAST_SEQ;
                    else if ((at_end == 1'b1))
                        reg_fstate <= BOT_SEQ;
                    else if ((pb_seq_up == 1'b1 && last_ram == 1'b1))
                        reg_fstate <= INIT;
                    else if ((at_end == 1'b0))
                        reg_fstate <= IN_SEQ;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= IN_SEQ;

                    addr_inc <= 1'b1;
                    at_end_rst <= 1'b0;
                    load <= 1'b0;
                end
                BOT_SEQ: begin
                    if ((at_end == 1'b0))
                        reg_fstate <= IN_SEQ;
                    else if ((pb_seq_up == 1'b1 && pb_seq_dn = 1'b0))
                        reg_fstate <= NEXT_SEQ;
                    else if ((pb_seq_dn == 1'b1 && pb_seq_up = 1'b0))
                        reg_fstate <= PREV_SEQ;
                    else if ((pb_seq_dn == 1'b1 && addr == 10'b00_0000_0000))
                        reg_fstate <= LAST_SEQ;
                    else if ((pb_seq_up == 1'b1 && last_ram == 1'b1))
                        reg_fstate <= INIT;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= BOT_SEQ;

                    at_end_rst <= 1'b1;
                    //addr <= start[9:0];

                    load <= 1'b1;
                end
                NEXT_SEQ: begin
                    if ((pb_up == 0))
                        reg_fstate <= IN_SEQ;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= NEXT_SEQ;

                    //addr <= start[9:0];

                    load <= 1'b1;
                    ram_counter_inc <= 1'b1;
					
					
                end
                PREV_SEQ: begin
                    if ((pb_seq_dn == 0))
                        reg_fstate <= IN_SEQ;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= PREV_SEQ;

                    ram_counter_dec <= 1'b1;

                    //addr <= start[9:0];

                    load <= 1'b1;
                end
                LAST_SEQ: begin
                    if ((pb_seq_dn == 0 && first_ram == 0))
                        reg_fstate <= IN_SEQ;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= LAST_SEQ;

                    ram_counter <= length[5:0];

                    addr <= start[9:0];

                    load <= 1'b1;
                end
                default: begin
                    load <= 1'bx;
                    addr <= 10'bxxxxxxxxxx;
                    ram_counter <= 6'bxxxxxx;
                    at_end_rst <= 1'bx;
                    addr_inc <= 1'bx;
                    ram_counter_inc <= 1'bx;
                    ram_counter_dec <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // ROM_state
